interface if_dut ();
    logic clk;
    logic rstn;
    logic in;
    logic out;
endinterface