interface if_dut (input clk);
    logic clk;
    logic rstn;
    logic in;
    logic out;
endinterface